LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY RCA4Bit IS
    PORT (
        Cin0:

        A0:
        A1:
        A2:
        A3:

        B0:
        B1:
        B2:
        B3:

    );

END RCA4Bit;
--
--
---------------------------------------
--
--
ARCHITECTURE Behaviour OF RCA4Bit IS
BEGIN

END Behaviour;