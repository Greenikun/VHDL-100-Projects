LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY NOT_GATE IS
    PORT (
        A : IN STD_LOGIC;
        Y : OUT STD_LOGIC
    );
END NOT_GATE;

ARCHITECTURE behavioural OF NOT_GATE IS
BEGIN
    Y <= NOT A;
END behavioural;