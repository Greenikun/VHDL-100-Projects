LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY FullAdder_tb IS
END FullAdder_tb;
--
--
----------------------------------------------------
--
--
ARCHITECTURE Test OF FullAdder_tb IS
BEGIN
END Test;